*DAC R-2R


***********OPAMP***********************
M1 2 2 1 1 pfet W=12U L=0.2u
M2 3 2 1 1  pfet W=12U L=0.2u
M3 2 out 6 1x nfet W=18U L=0.2u
M4 3 in_p 6 1x nfet W=18U L=0.2u
M5 6 7 1x 1x nfet W=1U L=1u
************NEEDS TO BE CHANGED
Rx1 1 7 2MEG
M7 7 7 1x 1x  nfet W=1U L=1u
M8 out 3 1 1 pfet W=20U L=0.2u
C1 3 out 2pf
M9 out 7 1x 1x nfet W=0.4U L=0.2u
Vdd 1 0 3.3V
************NEEDS TO BE CHANGED
Vss 1x 0 -3.3V
***********OPAMP***********************

R1 D9_ in_p 18k
R2 i in_p 9k
R3 D8_ i 18k
R4 h i 9k
R5 D7_ h 18k
R6 g h 9k
R7 D6_ g 18k
R8 f g 9k
R9 D5_ f 18k
R10 e f 9k
R11 D4_ e 18k
R12 d e 9k
R13 D3_ d 18k
R14 c d 9k
R15 D2_ c 18k
R16 b c 9k
R17 D1_ b 18k
R18 a b 9k
R19 D0_ a 18k
R20 a 0 18k

X1  D0 D0_ vref 1 0 switch
X2  D1 D1_ vref 1 0 switch
X3  D2 D2_ vref 1 0 switch
X4  D3 D3_ vref 1 0 switch
X5  D4 D4_ vref 1 0 switch
X6  D5 D5_ vref 1 0 switch
X7  D6 D6_ vref 1 0 switch
X8  D7 D7_ vref 1 0 switch
X9  D8 D8_ vref 1 0 switch
X10 D9 D9_ vref 1 0 switch

V9 D9 0 1.8V
V8 D8 0 1.8V
V7 D7 0 1.8V
V6 D6 0 1.8V
V5 D5 0 1.8V
V4 D4 0 1.8V
V3 D3 0 1.8V
V2 D2 0 1.8V
V1 D1 0 1.8V
V0 D0 0 1.8V

Vd_vref vref 0 3.3V
.SUBCKT switch data node vref s o
m1t node data_bar vref s pfet W=4u L=0.2u
m2t node data_bar o o nfet W=1u L=0.2u

m3t data_bar data s s pfet W=1.2u L=0.2u
m4t data_bar data o o nfet W=0.6u L=0.2u
.ENDS switch

.include osu018.lib
.tran 1ns 103us
.end