
*
.subckt DFFSR gnd vdd D S_ R_ Q CLK
Msp S S_ vdd vdd pfet w=2u l=0.2u
Msn S S_ gnd gnd nfet w=1u l=0.2u
Mrp R R_ vdd vdd pfet w=2u l=0.2u
Mrn R R_ gnd gnd nfet w=1u l=0.2u
M0 a_2_6# R vdd vdd pfet w=2u l=0.2u
M1 vdd a_10_61# a_2_6# vdd pfet w=2u l=0.2u
M2 a_10_61# a_23_27# vdd vdd pfet w=2u l=0.2u
M3 vdd S a_10_61# vdd pfet w=2u l=0.2u
M4 a_23_27# a_47_71# a_2_6# vdd pfet w=1u l=0.2u
M5 a_57_6# a_47_4# a_23_27# vdd pfet w=1u l=0.2u
M6 vdd D a_57_6# vdd pfet w=2u l=0.2u
M7 vdd a_47_71# a_47_4# vdd pfet w=2u l=0.2u
M8 a_47_71# CLK vdd vdd pfet w=2u l=0.2u
M9 a_105_6# a_47_71# a_10_61# vdd pfet w=1u l=0.2u
M10 a_113_6# a_47_4# a_105_6# vdd pfet w=1u l=0.2u
M11 a_122_6# a_105_6# vdd vdd pfet w=2u l=0.2u
M12 vdd R a_122_6# vdd pfet w=2u l=0.2u
M13 a_113_6# a_122_6# vdd vdd pfet w=2u l=0.2u
M14 vdd S a_113_6# vdd pfet w=2u l=0.2u
M15 vdd a_122_6# Q vdd pfet w=2u l=0.2u
M16 a_10_6# R a_2_6# gnd nfet w=2u l=0.2u
M17 gnd a_10_61# a_10_6# gnd nfet w=2u l=0.2u
M18 a_26_6# a_23_27# gnd gnd nfet w=2u l=0.2u
M19 a_10_61# S a_26_6# gnd nfet w=2u l=0.2u
M20 a_23_27# a_47_4# a_2_6# gnd nfet w=1u l=0.2u
M21 a_57_6# a_47_71# a_23_27# gnd nfet w=1u l=0.2u
M22 gnd D a_57_6# gnd nfet w=1u l=0.2u
M23 gnd a_47_71# a_47_4# gnd nfet w=1u l=0.2u
M24 a_47_71# CLK gnd gnd nfet w=1u l=0.2u
M25 a_105_6# a_47_4# a_10_61# gnd nfet w=1u l=0.2u
M26 a_113_6# a_47_71# a_105_6# gnd nfet w=1u l=0.2u
M27 a_130_6# a_105_6# a_122_6# gnd nfet w=2u l=0.2u
M28 gnd R a_130_6# gnd nfet w=2u l=0.2u
M29 a_146_6# a_122_6# gnd gnd nfet w=2u l=0.2u
M30 a_113_6# S a_146_6# gnd nfet w=2u l=0.2u
M31 gnd a_122_6# Q gnd nfet w=1u l=0.2u
.ends DFFSR
.tran 3us

.include osu018.lib
