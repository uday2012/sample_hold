*AND

X1 Vdd_d 0 v_a v_b OUT AND

.subckt AND N001 0 N003 N004 OUT
M1 N001 N003 N002 N001 pfet l=0.2u w=2u
M2 N001 N004 N002 N001 pfet l=0.2u w=2u
M3 N002 N003 N005 0 nfet l=0.2u w=1u
M5 N001 N002 OUT N001 pfet l=0.2u w=2u
M6 OUT N002 0 0 nfet l=0.2u w=1u

M4 N005 N004 0 0 nfet l=0.2u w=1u
.ends AND

Va v_a  0 PULSE(0 1.8v 1ns 1ns 1ns 0.25us 0.5us)
Vb v_b 0 1.8v
Vdd Vdd_d 0 1.8v

.tran 5us
.inc osu018.lib

.control
run
plot V(OUT) V(v_a) V(v_b)
.endc
.end
