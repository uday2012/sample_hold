*DAC R-2R


***********OPAMP***********************
M1 3 2 1 1 pfet W=54u L=0.2u
M2 4 in_n 3 1 pfet W=27u L=0.2u
M3 5 in_p 3 1 pfet W=27u L=0.2u
M4 4 4 0 0 nfet W=6.75u L=0.2u
M5 5 4 0 0 nfet W=6.75u L=0.2u
M6 6 2 1 1 pfet W=54u L=0.2u
M7 6 5 0 0 nfet W=13.2u L=0.2u
Rz 5 x 500
Cc x 6 2.7pF
M8 1 6 out 0 nfet W=10u L=0.2u
M9 out 8 0 0 nfet W=0.4u L=0.2u
M10 2 2 1 1 pfet W=9u L=0.2u
I1 1 9 50u
M11 9 9 8 0 nfet W=25u L=0.2u
M12 2 9 10 0 nfet W=25u L=0.2u
M13 8 8 0 0 nfet W=2.5u L=0.2u
M14 10 8 0 0 nfet W=2.5u L=0.2u
Rf in_n out 2k
Rx in_n 0 2K
***********OPAMP***********************
Vdd 1 0 3.3V
.param lmin=0.2u

R1 D9_ in_p 18k
R2 i in_p 9k
R3 D8_ i 18k
R4 h i 9k
R5 D7_ h 18k
R6 g h 9k
R7 D6_ g 18k
R8 f g 9k
R9 D5_ f 18k
R10 e f 9k
R11 D4_ e 18k
R12 d e 9k
R13 D3_ d 18k
R14 c d 9k
R15 D2_ c 18k
R16 b c 9k
R17 D1_ b 18k
R18 a b 9k
R19 D0_ a 18k
R20 a 0 18k

X1  D0 D0_ vref 1 0 switch
X2  D1 D1_ vref 1 0 switch
X3  D2 D2_ vref 1 0 switch
X4  D3 D3_ vref 1 0 switch
X5  D4 D4_ vref 1 0 switch
X6  D5 D5_ vref 1 0 switch
X7  D6 D6_ vref 1 0 switch
X8  D7 D7_ vref 1 0 switch
X9  D8 D8_ vref 1 0 switch
X10 D9 D9_ vref 1 0 switch

V9 D9 0 PULSE(1.8V 0 1p 1n 1n 51200n 102400n)
V8 D8 0 PULSE(1.8V 0 1p 1n 1n 25600n 51200n)
V7 D7 0 PULSE(1.8V 0 1p 1n 1n 12800n 25600n)
V6 D6 0 PULSE(1.8V 0 1p 1n 1n 6400n 12800n)
V5 D5 0 PULSE(1.8V 0 1p 1n 1n 3200n 6400n)
V4 D4 0 PULSE(1.8V 0 1p 1n 1n 1600n 3200n)
V3 D3 0 PULSE(1.8V 0 1p 1n 1n 800n 1600n)
V2 D2 0 PULSE(1.8V 0 1p 1n 1n 400n 800n)
V1 D1 0 PULSE(1.8V 0 1p 1n 1n 200n 400n)
V0 D0 0 PULSE(1.8V 0 1p 1n 1n 100n 200n)

Vd_vref vref 0 3.3V

.SUBCKT switch data node vref s o
m1t node data_bar vref s pfet W=4u L=0.2u
m2t node data_bar o o nfet W=1u L=0.2u

m3t data_bar data s s pfet W=1.2u L=0.2u
m4t data_bar data o o nfet W=0.6u L=0.2u
.ENDS switch

.include osu018.lib
.tran 1ns 20us
.end